module bpm_detection #(
    threshold = 
)