//module seven_segment_display #(
    
//)(

//);